`include "ha.sv"

module test (
	output wire [7:0] res [1:0],
	input wire [19:0] values [2:0]
);

	always @(values[0], values[1]) begin
		for(integer ;)
	end

endmodule
