/* Dadda Tree module
 * It performs the multioperand additions
 * in a CSA-style and provides two unsigned 
 * numbers for the final addition
 */

module dadda_tree (
	output reg [47:0] daddares [0:1],
	input wire [47:0] daddamat [0:8]
);
	
endmodule